module rotor();
endmodule