module EnigmaMachine();
endmodule

module rotor();
endmodule
