module EnigmaMachine();
endmodule